module test (
    input test
);
    
endmodule